`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:28:17 08/11/2021 
// Design Name: 
// Module Name:    ControlUnit 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ControlUnit( input [3:0]OpCode,
						  input [2:0]Function,
						  output reg [2:0] ALU,
						  output reg OUTLD, MWE, WE, S1,S2,S3,S4,S5,S6,S7,S8,S9 ); // s4	s5	s3	s2	s1	s9	WE	s6	s7	s8	ALU2	ALU1	ALU0	MWE	OUTLD
	
	always @(*)
	begin
		case (OpCode)
			4'b0000: 
			begin
				case (Function)
					3'b000: 
					begin
						S4=1;
						S5=0;
						S3=0;
						S2=0;
						S1=0;
						S9=0;
						WE=1;
						S6=0;
						S7=1;
						S8=0;
						ALU=3'b000;
						MWE=0;
						OUTLD=0;
					end
					3'b001:
					begin
						S4=1;
						S5=0;
						S3=0;
						S2=0;
						S1=0;
						S9=0;
						WE=1;
						S6=0;
						S7=1;
						S8=0;
						ALU=3'b001;
						MWE=0;
						OUTLD=0;
					end 
					3'b010: 
					begin 
						S4=1;
						S5=0;
						S3=0;
						S2=0;
						S1=0;
						S9=0;
						WE=1;
						S6=0;
						S7=1;
						S8=0;
						ALU=3'b010;
						MWE=0;
						OUTLD=0;
					end
					
					3'b011:
					begin
						S4=1;
						S5=0;
						S3=0;
						S2=0;
						S1=0;
						S9=0;
						WE=1;
						S6=0;
						S7=1;
						S8=0;
						ALU=3'b011;
						MWE=0;
						OUTLD=0;
					end

					3'b100: 
					begin
						S4=1;
						S5=0;
						S3=0;
						S2=0;
						S1=0;
						S9=0;
						WE=1;
						S6=0;
						S7=1;
						S8=0;
						ALU=3'b100;
						MWE=0;
						OUTLD=0;
					end
					3'b101: 
					begin
						S4=1;
						S5=0;
						S3=0;
						S2=0;
						S1=0;
						S9=0;
						WE=1;
						S6=0;
						S7=1;
						S8=0;
						ALU=3'b101;
						MWE=0;
						OUTLD=0;
					end
					3'b110: 
					begin
						S4=1;
						S5=0;
						S3=0;
						S2=0;
						S1=0;
						S9=0;
						WE=1;
						S6=0;
						S7=1;
						S8=0;
						ALU=3'b110;
						MWE=0;
						OUTLD=0;
					end
					3'b111: 
					begin
						S4=1;
						S5=0;
						S3=0;
						S2=0;
						S1=0;
						S9=0;
						WE=1;
						S6=0;
						S7=1;
						S8=0;
						ALU=3'b111;
						MWE=0;
						OUTLD=0;
					end
				endcase
			end
			4'b0100:
			begin
				S4=0;
				S5=0;
				S3=0;
				S2=0;
				S1=0;
				S9=0;
				WE=1;
				S6=0;
				S7=1;
				S8=1;
				ALU=3'b000;
				MWE=0;
				OUTLD=0;
			end
			4'b0101:
			begin
				S4=0;
				S5=0;
				S3=0;
				S2=0;
				S1=0;
				S9=0;
				WE=1;
				S6=0;
				S7=1;
				S8=1;
				ALU=3'b010;
				MWE=0;
				OUTLD=0;
			end
			4'b0110:
			begin
				S4=0;
				S5=0;
				S3=0;
				S2=0;
				S1=0;
				S9=0;
				WE=1;
				S6=0;
				S7=1;
				S8=1;
				ALU=3'b011;
				MWE=0;
				OUTLD=0;
			end
			4'b0111:
			begin
				S4=0;
				S5=0;
				S3=0;
				S2=0;
				S1=0;
				S9=0;
				WE=1;
				S6=0;
				S7=0;
				S8=1;
				ALU=3'b000;
				MWE=0;
				OUTLD=0;		
			end
			4'b1000:
			begin
				S4=0;
				S5=0;
				S3=0;
				S2=0;
				S1=0;
				S9=0;
				WE=0;
				S6=0;
				S7=0;
				S8=1;
				ALU=3'b000;
				MWE=1;
				OUTLD=0;
			end
			4'b1011:
			begin
				S4=0;
				S5=0;
				S3=0;
				S2=1;
				S1=0;
				S9=0;
				WE=0;
				S6=0;
				S7=0;
				S8=0;
				ALU=3'b000;
				MWE=0;
				OUTLD=0;
			end
			4'b1100:
			begin
				S4=0;
				S5=1;
				S3=0;
				S2=1;
				S1=0;
				S9=0;
				WE=1;
				S6=0;
				S7=0;
				S8=0;
				ALU=3'b000;
				MWE=0;
				OUTLD=0;
			end
			4'b0011:
			begin
				S4=0;
				S5=0;
				S3=0;
				S2=1;
				S1=1;
				S9=0;
				WE=0;
				S6=0;
				S7=0;
				S8=0;
				ALU=3'b000;
				MWE=0;
				OUTLD=0;
			end
			4'b1001:
			begin
				S4=0;
				S5=0;
				S3=0;
				S2=0;
				S1=1;
				S9=1;
				WE=0;
				S6=0;
				S7=0;
				S8=0;
				ALU=3'b001;
				MWE=0;
				OUTLD=0;
			end
			4'b1010:
			begin
				S4=0;
				S5=0;
				S3=0;
				S2=0;
				S1=1;
				S9=0;
				WE=0;
				S6=0;
				S7=0;
				S8=0;
				ALU=3'b001;
				MWE=0;
				OUTLD=0;
			end
			4'b0001:
			begin
				S4=1;
				S5=0;
				S3=0;
				S2=0;
				S1=0;
				S9=0;
				WE=1;
				S6=1;
				S7=1;
				S8=0;
				ALU=3'b000;
				MWE=0;
				OUTLD=0;
			end
			4'b0010:
			begin
				S4=0;
				S5=0;
				S3=0;
				S2=0;
				S1=0;
				S9=0;
				WE=0;
				S6=0;
				S7=0;
				S8=0;
				ALU=3'b000;
				MWE=0;
				OUTLD=1;
			end
			4'b1110:
			begin
				S4=0;
				S5=0;
				S3=0;
				S2=0;
				S1=0;
				S9=0;
				WE=0;
				S6=0;
				S7=0;
				S8=0;
				ALU=3'b000;
				MWE=0;
				OUTLD=0;
			end
			4'b1111:
			begin
				S4=0;
				S5=0;
				S3=1;
				S2=0;
				S1=0;
				S9=0;
				WE=0;
				S6=0;
				S7=0;
				S8=0;
				ALU=3'b000;
				MWE=0;
				OUTLD=0;
			end
			default:
			begin
				S4=0;
				S5=0;
				S3=0;
				S2=0;
				S1=0;
				S9=0;
				WE=0;
				S6=0;
				S7=0;
				S8=0;
				ALU=3'b000;
				MWE=0;
				OUTLD=0;
			end
			endcase
	end

endmodule
